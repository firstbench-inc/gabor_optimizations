  parameter  coeff1_int_mult1 = 2,
  parameter  coeff1_dec_mult1 = 15,
  parameter  coeff1_int_mult2 = 2,
  parameter  coeff1_dec_mult2 = 15,
  parameter  coeff1_int_mult3 = 2,
  parameter  coeff1_dec_mult3 = 15,
  parameter  coeff1_int_mult4 = 2,
  parameter  coeff1_dec_mult4 = 15,
  parameter  coeff1_int_mult5 = 2,
  parameter  coeff1_dec_mult5 = 15,
  parameter  coeff1_int_mult6 = 2,
  parameter  coeff1_dec_mult6 = 15,
  parameter  coeff1_int_mult7 = 2,
  parameter  coeff1_dec_mult7 = 15,
  parameter  coeff1_int_mult8 = 2,
  parameter  coeff1_dec_mult8 = 15,
  parameter  pixel_int_width = 9,
  parameter  pixel_dec_width = 0,
  parameter  col_adder_width = 22

//  parameter  coeff1_int_mult9 = 2,
 // parameter  coeff1_dec_mult9 = 15,
  //parameter  coeff1_int_mult10 = 2,
  //parameter  coeff1_dec_mult10 = 15,
  //parameter  coeff1_int_mult11 = 2,
  //parameter  coeff1_dec_mult11 = 15,
  //parameter  coeff1_int_mult12 = 2,
  //parameter  coeff1_dec_mult12 = 15,
  //parameter  coeff1_int_mult13 = 2,
  //parameter  coeff1_dec_mult13 = 15,
// parameter ex
