module lut();
endmodule
